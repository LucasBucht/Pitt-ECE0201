--
-- VHDL Entity CPU_Design_lib.FiveBitCounter.arch_name
--
-- Created:
--          by - lmb290.UNKNOWN (SSOE-COELABS17)
--          at - 14:36:25 12/ 8/2025
--
-- using Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 17:42:50
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY FiveBitCounter IS
   PORT( 
      clock : IN     std_logic;
      reset : IN     std_logic;
      count : OUT    std_logic_vector (4 DOWNTO 0)
   );

-- Declarations

END FiveBitCounter ;


--
-- VHDL Architecture CPU_Design_lib.FiveBitCounter.fsm
--
-- Created:
--          by - lmb290.UNKNOWN (SSOE-COELABS17)
--          at - 15:24:44 12/ 8/2025
--
-- Generated by Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 17:42:50
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
 
ARCHITECTURE fsm OF FiveBitCounter IS

   TYPE STATE_TYPE IS (
      s0,
      s1,
      s2,
      s3,
      s4,
      s5,
      s6,
      s7,
      s8,
      s9,
      s10,
      s11,
      s12,
      s13,
      s14,
      s15,
      s16,
      s17,
      s18,
      s19,
      s20
   );
 
   -- Declare current and next state signals
   SIGNAL current_state : STATE_TYPE;
   SIGNAL next_state : STATE_TYPE;

BEGIN

   -----------------------------------------------------------------
   clocked_proc : PROCESS ( 
      clock,
      reset
   )
   -----------------------------------------------------------------
   BEGIN
      IF (reset = '0') THEN
         current_state <= s0;
      ELSIF (clock'EVENT AND clock = '1') THEN
         current_state <= next_state;
      END IF;
   END PROCESS clocked_proc;
 
   -----------------------------------------------------------------
   nextstate_proc : PROCESS ( 
      current_state
   )
   -----------------------------------------------------------------
   BEGIN
      CASE current_state IS
         WHEN s0 => 
            next_state <= s1;
         WHEN s1 => 
            next_state <= s2;
         WHEN s2 => 
            next_state <= s3;
         WHEN s3 => 
            next_state <= s4;
         WHEN s4 => 
            next_state <= s5;
         WHEN s5 => 
            next_state <= s6;
         WHEN s6 => 
            next_state <= s7;
         WHEN s7 => 
            next_state <= s8;
         WHEN s8 => 
            next_state <= s9;
         WHEN s9 => 
            next_state <= s10;
         WHEN s10 => 
            next_state <= s11;
         WHEN s11 => 
            next_state <= s12;
         WHEN s12 => 
            next_state <= s13;
         WHEN s13 => 
            next_state <= s14;
         WHEN s14 => 
            next_state <= s15;
         WHEN s15 => 
            next_state <= s16;
         WHEN s16 => 
            next_state <= s17;
         WHEN s17 => 
            next_state <= s18;
         WHEN s18 => 
            next_state <= s19;
         WHEN s19 => 
            next_state <= s20;
         WHEN s20 => 
            next_state <= s0;
         WHEN OTHERS =>
            next_state <= s0;
      END CASE;
   END PROCESS nextstate_proc;
 
   -----------------------------------------------------------------
   output_proc : PROCESS ( 
      current_state
   )
   -----------------------------------------------------------------
   BEGIN

      -- Combined Actions
      CASE current_state IS
         WHEN s0 => 
            count <= "00000";
         WHEN s1 => 
            count <= "00001";
         WHEN s2 => 
            count <= "00010";
         WHEN s3 => 
            count <= "00011";
         WHEN s4 => 
            count <= "00100";
         WHEN s5 => 
            count <= "00101";
         WHEN s6 => 
            count <= "00110";
         WHEN s7 => 
            count <= "00111";
         WHEN s8 => 
            count <= "01000";
         WHEN s9 => 
            count <= "01001";
         WHEN s10 => 
            count <= "01010";
         WHEN s11 => 
            count <= "01011";
         WHEN s12 => 
            count <= "01100";
         WHEN s13 => 
            count <= "01101";
         WHEN s14 => 
            count <= "01110";
         WHEN s15 => 
            count <= "01111";
         WHEN s16 => 
            count <= "10000";
         WHEN s17 => 
            count <= "10001";
         WHEN s18 => 
            count <= "10010";
         WHEN s19 => 
            count <= "10011";
         WHEN s20 => 
            count <= "10100";
         WHEN OTHERS =>
            NULL;
      END CASE;
   END PROCESS output_proc;
 
END fsm;
