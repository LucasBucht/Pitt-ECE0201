--
-- VHDL Entity CPU_Design_lib.FSM_Controller.arch_name
--
-- Created:
--          by - lmb290.UNKNOWN (SSOE-COELABS19)
--          at - 13:18:58 11/20/2025
--
-- using Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 17:42:50
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY FSM_Controller IS
   PORT( 
      clk           : IN     std_logic;
      data_in       : IN     std_logic_vector (8 DOWNTO 0);
      en            : IN     std_logic;
      rst           : IN     std_logic;
      ALU_Op        : OUT    std_logic_vector (2 DOWNTO 0);
      A_en          : OUT    std_logic;
      Bus_Sel       : OUT    std_logic_vector (1 DOWNTO 0);
      F_en          : OUT    std_logic;
      IR_en         : OUT    std_logic;
      Read_Address  : OUT    std_logic_vector (2 DOWNTO 0);
      Write_Address : OUT    std_logic_vector (2 DOWNTO 0);
      done          : OUT    std_logic
   );

-- Declarations

END FSM_Controller ;


--
-- VHDL Architecture CPU_Design_lib.FSM_Controller.fsm
--
-- Created:
--          by - lmb290.UNKNOWN (SSOE-COELABS19)
--          at - 14:24:50 12/ 4/2025
--
-- Generated by Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 17:42:50
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
 
ARCHITECTURE fsm OF FSM_Controller IS

   TYPE STATE_TYPE IS (
      Fetch,
      mvi,
      mv,
      ALU_A,
      Add,
      Sub,
      And_Op,
      Or_Op,
      Inv_Op,
      WriteBack
   );
 
   -- Declare current and next state signals
   SIGNAL current_state : STATE_TYPE;
   SIGNAL next_state : STATE_TYPE;

BEGIN

   -----------------------------------------------------------------
   clocked_proc : PROCESS ( 
      clk,
      rst
   )
   -----------------------------------------------------------------
   BEGIN
      IF (rst = '1') THEN
         current_state <= Fetch;
      ELSIF (clk'EVENT AND clk = '0') THEN
         IF (en = '1') THEN
            current_state <= next_state;
         END IF;
      END IF;
   END PROCESS clocked_proc;
 
   -----------------------------------------------------------------
   nextstate_proc : PROCESS ( 
      current_state,
      data_in,
      en
   )
   -----------------------------------------------------------------
   BEGIN
      CASE current_state IS
         WHEN Fetch => 
            IF ((data_in (8 downto 6) = "001") AND (en = '1')) THEN 
               next_state <= mvi;
            ELSIF ((data_in (8 downto 6) = "000") AND (en = '1')) THEN 
               next_state <= mv;
            ELSIF ((en = '1') AND NOT (data_in (8 downto 6) = "000") AND NOT (data_in (8 downto 6) = "001")) THEN 
               next_state <= ALU_A;
            ELSE
               next_state <= Fetch;
            END IF;
         WHEN mvi => 
            next_state <= Fetch;
         WHEN mv => 
            next_state <= Fetch;
         WHEN ALU_A => 
            IF ((en = '1') AND (data_in (8 downto 6) = "010")) THEN 
               next_state <= Add;
            ELSIF ((en = '1') AND (data_in (8 downto 6) = "011")) THEN 
               next_state <= Sub;
            ELSIF ((en = '1') AND (data_in (8 downto 6) = "110")) THEN 
               next_state <= And_Op;
            ELSIF ((en = '1') AND (data_in (8 downto 6) = "100")) THEN 
               next_state <= Or_Op;
            ELSIF ((en = '1') AND (data_in (8 downto 6) = "101")) THEN 
               next_state <= Inv_Op;
            ELSE
               next_state <= ALU_A;
            END IF;
         WHEN Add => 
            next_state <= WriteBack;
         WHEN Sub => 
            next_state <= WriteBack;
         WHEN And_Op => 
            next_state <= WriteBack;
         WHEN Or_Op => 
            next_state <= WriteBack;
         WHEN Inv_Op => 
            next_state <= WriteBack;
         WHEN WriteBack => 
            next_state <= Fetch;
         WHEN OTHERS =>
            next_state <= Fetch;
      END CASE;
   END PROCESS nextstate_proc;
 
   -----------------------------------------------------------------
   output_proc : PROCESS ( 
      current_state,
      data_in
   )
   -----------------------------------------------------------------
   BEGIN

      -- Combined Actions
      CASE current_state IS
         WHEN Fetch => 
            ALU_Op <= "000";
            F_en <= '0';
            Bus_Sel  <= "01";
            IR_en <=  '1';
            A_en <= '0';
            Read_Address <= "000";
            Write_Address <= "000";
            done <= '0';
         WHEN mvi => 
            ALU_Op <= "000";
            F_en <= '0';
            Bus_Sel  <= "01";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= "000";
            Write_Address <= data_in (5 downto 3);
            done <= '1';
         WHEN mv => 
            ALU_Op <= "000";
            F_en <= '0';
            Bus_Sel  <= "10";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= data_in (2 downto 0);
            Write_Address <= data_in (5 downto 3);
            done <= '1';
         WHEN ALU_A => 
            ALU_Op <= "000";
            F_en <= '0';
            Bus_Sel  <= "10";
            IR_en <=  '0';
            A_en <= '1';
            Read_Address <= data_in (5 downto 3);
            Write_Address <= data_in (5 downto 3);
            done <= '0';
         WHEN Add => 
            ALU_Op <= "000";
            F_en <= '1';
            Bus_Sel  <= "01";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= data_in(2 downto 0);
            Write_Address <= data_in(2 downto 0);
            done <= '0';
         WHEN Sub => 
            ALU_Op <= "100";
            F_en <= '1';
            Bus_Sel  <= "01";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= data_in(2 downto 0);
            Write_Address <= data_in(2 downto 0);
            done <= '0';
         WHEN And_Op => 
            ALU_Op <= "001";
            F_en <= '1';
            Bus_Sel  <= "01";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= data_in(2 downto 0);
            Write_Address <= data_in(2 downto 0);
            done <= '0';
         WHEN Or_Op => 
            ALU_Op <= "010";
            F_en <= '1';
            Bus_Sel  <= "01";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= data_in(2 downto 0);
            Write_Address <= data_in(2 downto 0);
            done <= '0';
         WHEN Inv_Op => 
            ALU_Op <= "011";
            F_en <= '1';
            Bus_Sel  <= "01";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= data_in(2 downto 0);
            Write_Address <= data_in(2 downto 0);
            done <= '0';
         WHEN WriteBack => 
            ALU_Op <= "000";
            F_en <= '0';
            Bus_Sel  <= "00";
            IR_en <=  '0';
            A_en <= '0';
            Read_Address <= "000";
            Write_Address <= data_in(5 downto 3);
            done <= '1';
         WHEN OTHERS =>
            NULL;
      END CASE;
   END PROCESS output_proc;
 
END fsm;
