--
-- VHDL Entity CPU_Design_lib.FSM_Controller.arch_name
--
-- Created:
--          by - lmb290.UNKNOWN (SSOE-COELABS19)
--          at - 13:18:58 11/20/2025
--
-- using Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 17:42:50
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY FSM_Controller IS
   PORT( 
      clk           : IN     std_logic;
      data_in       : IN     std_logic_vector (8 DOWNTO 0);
      en            : IN     std_logic;
      rst           : IN     std_logic;
      ALU_Op        : OUT    std_logic_vector (1 DOWNTO 0);
      A_en          : OUT    std_logic;
      Bus_Sel       : OUT    std_logic_vector (1 DOWNTO 0);
      F_en          : OUT    std_logic;
      IR_en         : OUT    std_logic;
      Read_Address  : OUT    std_logic_vector (2 DOWNTO 0);
      Write_Address : OUT    std_logic_vector (2 DOWNTO 0);
      done          : OUT    std_logic
   );

-- Declarations

END FSM_Controller ;


--
-- VHDL Architecture CPU_Design_lib.FSM_Controller.fsm
--
-- Created:
--          by - lmb290.UNKNOWN (SSOE-COELABS19)
--          at - 14:29:38 11/20/2025
--
-- Generated by Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 17:42:50
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;
 
ARCHITECTURE fsm OF FSM_Controller IS

   TYPE STATE_TYPE IS (
      Fetch,
      mvi
   );
 
   -- Declare current and next state signals
   SIGNAL current_state : STATE_TYPE;
   SIGNAL next_state : STATE_TYPE;

BEGIN

   -----------------------------------------------------------------
   clocked_proc : PROCESS ( 
      clk,
      rst
   )
   -----------------------------------------------------------------
   BEGIN
      IF (rst = '1') THEN
         current_state <= Fetch;
      ELSIF (clk'EVENT AND clk = '1') THEN
         IF (en = '1') THEN
            current_state <= next_state;
         END IF;
      END IF;
   END PROCESS clocked_proc;
 
   -----------------------------------------------------------------
   nextstate_proc : PROCESS ( 
      current_state,
      data_in
   )
   -----------------------------------------------------------------
   BEGIN
      CASE current_state IS
         WHEN Fetch => 
            IF (data_in (8 downto 6) = "001") THEN 
               next_state <= mvi;
            ELSE
               next_state <= Fetch;
            END IF;
         WHEN mvi => 
            next_state <= Fetch;
         WHEN OTHERS =>
            next_state <= Fetch;
      END CASE;
   END PROCESS nextstate_proc;
 
   -----------------------------------------------------------------
   output_proc : PROCESS ( 
      current_state,
      data_in
   )
   -----------------------------------------------------------------
   BEGIN

      -- Combined Actions
      CASE current_state IS
         WHEN Fetch => 
            IR_en <= '1';
            A_en <= '0';
            F_en <= '0';
            Done <= '0';
            Write_Address <= Data_In (5 downto 3);
         WHEN mvi => 
            IR_en <= '0';
            Bus_Sel <= "01";
            Done <= '1';
         WHEN OTHERS =>
            NULL;
      END CASE;
   END PROCESS output_proc;
 
END fsm;
