--
-- VHDL Entity CPU_Design_lib.FSM_Controller.arch_name
--
-- Created:
--          by - lmb290.UNKNOWN (SSOE-COELABS19)
--          at - 13:18:58 11/20/2025
--
-- using Siemens HDL Designer(TM) 2024.1 Built on 24 Jan 2024 at 17:42:50
--
LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.std_logic_arith.all;

ENTITY FSM_Controller IS
   PORT( 
      clk           : IN     std_logic;
      data_in       : IN     std_logic_vector (8 DOWNTO 0);
      en            : IN     std_logic;
      rst           : IN     std_logic;
      ALU_Op        : OUT    std_logic_vector (2 DOWNTO 0);
      A_en          : OUT    std_logic;
      Bus_Sel       : OUT    std_logic_vector (1 DOWNTO 0);
      F_en          : OUT    std_logic;
      IR_en         : OUT    std_logic;
      Read_Address  : OUT    std_logic_vector (2 DOWNTO 0);
      Write_Address : OUT    std_logic_vector (2 DOWNTO 0);
      Write_Enable  : OUT    std_logic;
      done          : OUT    std_logic
   );

-- Declarations

END FSM_Controller ;

